library verilog;
use verilog.vl_types.all;
entity SumV2_vlg_vec_tst is
end SumV2_vlg_vec_tst;
