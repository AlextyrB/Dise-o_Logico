library verilog;
use verilog.vl_types.all;
entity Multiplicador_vlg_vec_tst is
end Multiplicador_vlg_vec_tst;
